module OR(A, B, result);
    input [31:0] A, B;
    output [31:0] result;

    or OR0(result[0], A[0], B[0]);
    or OR1(result[1], A[1], B[1]);
    or OR2(result[2], A[2], B[2]);
    or OR3(result[3], A[3], B[3]);
    or OR4(result[4], A[4], B[4]);
    or OR5(result[5], A[5], B[5]);
    or OR6(result[6], A[6], B[6]);
    or OR7(result[7], A[7], B[7]);
    or OR8(result[8], A[8], B[8]);
    or OR9(result[9], A[9], B[9]);
    or OR10(result[10], A[10], B[10]);
    or OR11(result[11], A[11], B[11]);
    or OR12(result[12], A[12], B[12]);
    or OR13(result[13], A[13], B[13]);
    or OR14(result[14], A[14], B[14]);
    or OR15(result[15], A[15], B[15]);
    or OR16(result[16], A[16], B[16]);
    or OR17(result[17], A[17], B[17]);
    or OR18(result[18], A[18], B[18]);
    or OR19(result[19], A[19], B[19]);
    or OR20(result[20], A[20], B[20]);
    or OR21(result[21], A[21], B[21]);
    or OR22(result[22], A[22], B[22]);
    or OR23(result[23], A[23], B[23]);
    or OR24(result[24], A[24], B[24]);
    or OR25(result[25], A[25], B[25]);
    or OR26(result[26], A[26], B[26]);
    or OR27(result[27], A[27], B[27]);
    or OR28(result[28], A[28], B[28]);
    or OR29(result[29], A[29], B[29]);
    or OR30(result[30], A[30], B[30]);
    or OR31(result[31], A[31], B[31]);
endmodule