module AND(A, B, result);
    input [31:0] A, B;
    output [31:0] result;

    and AND0(result[0], A[0], B[0]);
    and AND1(result[1], A[1], B[1]);
    and AND2(result[2], A[2], B[2]);
    and AND3(result[3], A[3], B[3]);
    and AND4(result[4], A[4], B[4]);
    and AND5(result[5], A[5], B[5]);
    and AND6(result[6], A[6], B[6]);
    and AND7(result[7], A[7], B[7]);
    and AND8(result[8], A[8], B[8]);
    and AND9(result[9], A[9], B[9]);
    and AND10(result[10], A[10], B[10]);
    and AND11(result[11], A[11], B[11]);
    and AND12(result[12], A[12], B[12]);
    and AND13(result[13], A[13], B[13]);
    and AND14(result[14], A[14], B[14]);
    and AND15(result[15], A[15], B[15]);
    and AND16(result[16], A[16], B[16]);
    and AND17(result[17], A[17], B[17]);
    and AND18(result[18], A[18], B[18]);
    and AND19(result[19], A[19], B[19]);
    and AND20(result[20], A[20], B[20]);
    and AND21(result[21], A[21], B[21]);
    and AND22(result[22], A[22], B[22]);
    and AND23(result[23], A[23], B[23]);
    and AND24(result[24], A[24], B[24]);
    and AND25(result[25], A[25], B[25]);
    and AND26(result[26], A[26], B[26]);
    and AND27(result[27], A[27], B[27]);
    and AND28(result[28], A[28], B[28]);
    and AND29(result[29], A[29], B[29]);
    and AND30(result[30], A[30], B[30]);
    and AND31(result[31], A[31], B[31]);
endmodule