module SRA1_mult(A, result);
    input [64:0] A;
    output [64:0] result;

    assign result[64] = A[64];
    assign result[63] = A[64];
    assign result[62] = A[63];
    assign result[61] = A[62];
    assign result[60] = A[61];
    assign result[59] = A[60];
    assign result[58] = A[59];
    assign result[57] = A[58];
    assign result[56] = A[57];
    assign result[55] = A[56];
    assign result[54] = A[55];
    assign result[53] = A[54];
    assign result[52] = A[53];
    assign result[51] = A[52];
    assign result[50] = A[51];
    assign result[49] = A[50];
    assign result[48] = A[49];
    assign result[47] = A[48];
    assign result[46] = A[47];
    assign result[45] = A[46];
    assign result[44] = A[45];
    assign result[43] = A[44];
    assign result[42] = A[43];
    assign result[41] = A[42];
    assign result[40] = A[41];
    assign result[39] = A[40];
    assign result[38] = A[39];
    assign result[37] = A[38];
    assign result[36] = A[37];
    assign result[35] = A[36];
    assign result[34] = A[35];
    assign result[33] = A[34];
    assign result[32] = A[33];
    assign result[31] = A[32];
    assign result[30] = A[31];
    assign result[29] = A[30];
    assign result[28] = A[29];
    assign result[27] = A[28];
    assign result[26] = A[27];
    assign result[25] = A[26];
    assign result[24] = A[25];
    assign result[23] = A[24];
    assign result[22] = A[23];
    assign result[21] = A[22];
    assign result[20] = A[21];
    assign result[19] = A[20];
    assign result[18] = A[19];
    assign result[17] = A[18];
    assign result[16] = A[17];
    assign result[15] = A[16];
    assign result[14] = A[15];
    assign result[13] = A[14];
    assign result[12] = A[13];
    assign result[11] = A[12];
    assign result[10] = A[11];
    assign result[9] = A[10];
    assign result[8] = A[9];
    assign result[7] = A[8];
    assign result[6] = A[7];
    assign result[5] = A[6];
    assign result[4] = A[5];
    assign result[3] = A[4];
    assign result[2] = A[3];
    assign result[1] = A[2];
    assign result[0] = A[1];
endmodule