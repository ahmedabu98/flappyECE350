module isCollided(x